library verilog;
use verilog.vl_types.all;
entity VGA_Basis_v0_vlg_tst is
end VGA_Basis_v0_vlg_tst;
